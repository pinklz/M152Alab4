`timescale 1ns / 1ps

module ball(

    );
endmodule