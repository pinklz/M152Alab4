`timescale 1ns / 1ps

module clock_divider(

    );
endmodule