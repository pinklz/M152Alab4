`timescale 1ns / 1ps

module ball(
    input wire clk,
    input wire x_initial,
    input wire y_initial,
    input wire vx,
    input wire vy,

    output wire x_out,
    output wire y_out,
    );


endmodule