`timescale 1ns / 1ps

module board(

    );
endmodule