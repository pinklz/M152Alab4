`timescale 1ns / 1ps

module debouncer(

    );
endmodule