`timescale 1ns / 1ps

module physics_controller(
    
    );
endmodule